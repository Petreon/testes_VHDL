entity MUX2X1 is
	port (A: in bit; B: in bit; C: in bit; S: out bit);
end MUX2X1;