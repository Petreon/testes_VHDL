entity mux2x1 is
port (A,B,C: in bit; S: out bit);
end mux2x1;
