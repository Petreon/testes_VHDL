architecture algoritmica of dec4x16vetor is

begin
	process(E)
	begin
		case E is
		when "0000" => S <= "0000000000000001";
		when "0001" => S <= "0000000000000010";
		when "0010" => S <= "0000000000000100";
		when "0011" => S <= "0000000000001000";
		when "0100" => S <= "0000000000010000";
		when "0101" => S <= "0000000000100000";
		when "0110" => S <= "0000000001000000";
		when "0111" => S <= "0000000010000000";
		when "1000" => S <= "0000000100000000";
		when "1001" => S <= "0000001000000000";
		when "1010" => S <= "0000010000000000";
		when "1011" => S <= "0000100000000000";
		when "1100" => S <= "0001000000000000";
		when "1101" => S <= "0010000000000000";
		when "1110" => S <= "0100000000000000";
		when "1111" => S <= "1000000000000000";
		end case;
	end process;
end algoritmica;